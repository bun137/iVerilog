module basic_not(a, y);  
input a;
output y;
assign y = ! a;
endmodule
